module add_sub_1digit (result,c_out,sign,a,b,m,cin);
  input [4:0]a,b;
  input m,cin;
  output c_out,sign;
  output [3:0]result;
  wire [3:0]acomp,bcomp,s,s1,s3;
  wire t1,t2,t3,t4,ta,tb,Cout,s2,Cout1,Cout2,t5,t6,Cout3,t7,t8,t9,t10,t11,Cout4,L,E,G,t12,t13,t14,t_0,t_1,t_2,t_3;
  nor g1 (t1,0,a[4]);
  xor g2 (t2,b[4],m);
  nor g3 (ta,t1,t2);
  nines_complement g4 (a[3:0],ta,acomp);
  nor g5 (t3,t2,0);
  nor g6 (tb,t3,a[4]);
  nines_complement g7 (b[3:0],tb,bcomp);
  fulladd4 g8 (s,Cout,acomp,bcomp,cin);
  xor g9 (t4,ta,tb);
  fulladd4 g30 (s1,Cout1,s,({1'b0,t4,t4,t4}),1'b0);
  FAdd g31 (Cout,t4,Cout1,s2,Cout2);
  not g10 (t5,t4);
  nor g11 (t6,Cout2,t5);
  xor g12 (t_0,s1[0],t6);
  xor g13 (t_1,s1[1],t6);
  xor g14 (t_2,s1[2],t6);
  xor g15 (t_3,s1[3],t6);
  fulladd4 g16 (s3,Cout3,(4'b0000),({t_3,t_2,t_1,t_0}),t6);
  nand g17 (t7,s3[1],s3[3]);
  nand g18 (t8,s3[2],s3[3]);
  nand g19 (t9,t5,Cout);
  nand g20 (t10,t7,t8,t9);
  fulladd4 g21 (result,Cout4,s3,({1'b0,t10,t10,1'b0}),1'b0);
  not g22 (t11,Cout4);
  nand g23 (c_out,t11,t9);
  comparator_struct g24 (a[3:0],b[3:0],L,E,G);
  nand g25 (t12,L,t2);
  nand g26 (t13,a[4],G);
  nand g27 (t14,a[4],t2);
  nand g28 (sign,t12,t13,t14);
endmodule